﻿;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      27
619734.2,4239063.4,HWB
624348.3,4243212.4,SUT
615180.4,4216618.4,SLTRM004
624476.9,4208582.2,HOL
636491.6,4185281.5,ROLD059
614797.6,4223035.8,RSAC101
616952.5,4212848.6,FAL
625222.5,4203213.9,ROLD024
623598.2,4238356.2,SSS
636454.1,4186988.1,CHGRL009
629727.3,4233179.3,Georg_SL
629291.6,4192502.2,CHVCT000
615029,4212420.9,RSAN018
625718.9,4194688.9,ROLD034
630802.2,4234030.6,CHDCC000
647500.8,4192114.6,RSAN072
635762.3,4206110.6,TRN
618521.7,4214201.8,FCT
629664.2,4235427.1,RSAC128
630762.5,4257477,RSAC155
643575.2,4202944.9,RSAN058
629219.1,4233351.8,RSAC123
616676.6,4208098.2,SLDUT007
625274.8,4218552.5,MOK
639778,4185041,PDC
647096.2,4185827.7,ROLD074
597451.6,4219938,SLMZU025
