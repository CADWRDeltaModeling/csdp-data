;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      461
652291.3125,4172465.0,1
652401.1875000001,4174797.25,2
651800.6875,4176016.25,3
650044.0,4176792.75,4
649423.0,4179715.75,5
649669.1874999999,4182589.25,6
648443.8125,4184173.5,7
647237.0625,4185855.5,8
648354.25,4187713.0,9
647489.8125,4190138.5,10
647526.5,4192087.4999999995,11
646971.1875,4195317.5,12
647722.9375,4198306.0,13
646960.6875,4199204.5,14
646258.6875,4200263.0,15
645341.875,4200690.0,16
653984.1249999999,4170361.25,17
646236.5625,4201770.0,18
645129.75,4202089.5,19
644123.0,4202518.5,20
643233.6875,4203385.0,21
641995.25,4204667.5,22
640357.0,4205866.0,23
639403.5,4206340.0,24
637535.8125,4206248.5,25
636600.6875,4206649.0,26
636786.6875,4207985.0,27
635170.4375,4207343.5,28
635314.5625,4208409.5,29
634127.9375,4209928.5,30
632414.8125,4210196.0,31
632632.1875,4210997.5,32
631497.375,4211860.5,33
630043.0,4212840.0,34
628593.4375,4213038.5,35
628660.3125,4214299.5,36
627151.75,4213231.0,37
625286.5,4215502.5,38
625108.4375,4216137.5,39
624931.6875,4217185.5,40
621470.0,4218234.0,41
618784.375,4216400.5,42
615728.9375,4216061.0,43
615841.0625,4213249.5,44
611401.1875,4209956.0,45
604438.5,4208698.0,46
602633.0,4209643.5,47
646515.5000000001,4186410.5,48
646028.0625,4187282.5000000005,49
645366.375,4187263.5,50
644353.8125,4186947.75,51
643018.9375,4187291.75,52
642598.8125,4186989.5,53
641645.8125,4185910.75,54
640142.5,4185524.75,55
639159.9375,4186107.25,56
638985.6929687959,4185072.082274425,57
638937.5625,4184888.7500000005,58
637840.25,4184496.5,59
637057.6875,4184976.75,60
635696.5625,4184959.0000000005,61
634820.3125,4184459.75,62
634158.9375,4183453.7500000005,63
633404.9375,4182730.7499999995,64
632312.625,4182652.25,65
630772.125,4183653.5,66
629818.875,4184470.0,67
629153.5625,4185159.0,68
628267.0,4185764.0,69
626906.0625,4186453.0,70
627388.0625,4187144.5,71
627296.5625,4187984.0,72
627018.25,4188880.0,73
626758.3125,4189671.75,74
626353.3125,4190704.5,75
613113.8125,4208441.0,76
625478.4375,4191891.0,77
625077.6875,4193038.25,78
625216.5,4194337.5,79
626002.3125,4195060.5,80
625478.4375,4196111.0,81
626290.5,4197130.0,82
626916.5,4198102.0,84
626762.0,4199155.0,85
626466.0,4200158.0,86
626033.75,4200540.5,88
626058.5625,4201644.5,89
625184.3125,4201804.0,90
626087.6875,4202299.0,91
625435.375,4202776.5,92
625067.75,4203805.5,93
624563.1875,4204863.0,94
624716.25,4206435.5,97
625748.0,4207048.5,98
624676.5625,4207441.5,99
626698.8125,4208604.5,100
624976.5625,4211592.5,101
624560.75,4210245.5,102
624402.3125,4213537.5,103
642063.125,4188028.5,104
642572.5,4190194.0,105
642842.6875,4191531.2500000005,106
642203.75,4193334.25,107
641032.8125,4194434.5,108
639317.0625,4194633.5,109
637810.875,4195042.5,110
636603.3125,4194293.0,111
634764.4375,4193850.5,112
632826.0625,4194573.5,113
632289.0625,4195569.0,114
632118.8125,4196189.5,115
631128.625,4196582.5,116
630402.1875,4197315.0,117
630319.1875,4198020.5,118
629197.9375,4198380.5,119
629415.5,4199343.5,120
628896.875,4200205.0,121
628750.125,4201012.0,122
629630.3125,4201124.5,123
629145.6875,4202177.5,124
628739.6875,4203437.5,125
628642.75,4204614.0,126
628734.4375,4205384.0,127
629111.625,4206306.0,128
629837.25,4207034.0,129
630653.6875,4207075.5,130
630892.875,4207914.5,131
630164.6875,4208029.5,132
630122.75,4209242.5,133
629163.1875,4211556.5,134
630444.9375,4204553.5,135
630562.1875,4205460.5,136
631170.5625,4206185.5,137
643021.0,4200931.0,138
642342.5625,4202413.5,139
635471.6875,4205858.0,140
634030.875,4205002.5,141
633934.0625,4203728.5,142
632388.5625,4203731.0,143
630845.625,4203727.5,144
629680.0625,4203699.5,145
637839.6875,4199765.0,146
635919.625,4201887.0,147
634442.25,4202832.5,148
639074.3125,4183841.0000000005,149
639192.8125,4181795.25,150
645250.375,4181255.5,151
644446.375,4181696.75,152
643951.0,4181192.5,153
642975.375,4181314.0,154
642208.625,4181533.4999999995,155
641932.25,4182303.0,156
641365.7499999999,4181880.5,157
640666.625,4182830.75,158
640021.4375,4182442.5,159
639571.8125000001,4183094.5,160
648865.5,4180466.5,162
646494.0822180585,4182451.1615983737,163
645370.6875,4183844.0,164
643561.9284385688,4185100.083037729,165
645553.7373738948,4183113.321092806,166
643434.875,4184954.75,167
641475.5,4185418.25,168
639560.6875000001,4185177.25,169
640380.5625000001,4187039.75,170
638224.75,4186992.75,171
636503.75,4186942.75,172
635427.1875,4186922.0,173
634353.1875,4186903.5,174
633232.0625,4186877.5,175
632155.4375,4186851.25,176
630882.375,4186830.25,177
628810.375,4186798.75,178
625459.9375,4186288.75,179
624569.9375,4184215.7500000005,181
628383.4375,4188606.25,182
628737.0625,4189541.4999999995,183
628940.75,4190098.75,184
628333.6875,4190196.25,185
628358.5,4190951.75,186
627710.25,4190720.25,187
631754.6875,4193963.0,188
630458.0625,4193245.25,189
629606.75,4192766.0000000005,190
628783.3125,4192321.7500000005,191
627285.875,4191424.75,192
628936.125,4197245.0,194
627471.875,4197221.5,195
625049.875,4197728.5,196
623964.9375,4198022.5,197
622519.125,4197569.5,198
622319.625,4198858.5,199
622129.0625,4200201.0,200
622315.125,4201635.5,201
622667.0625,4202774.5,202
623460.5625,4203630.5,203
622512.375,4204128.5,204
621015.0,4204108.0,205
619354.0,4204025.0,206
628669.375,4207349.5,207
627032.6875,4207898.5,208
622959.5625,4188789.5,209
623872.6875,4189198.25,210
624501.375,4190044.25,211
624917.875,4191343.5000000005,212
627652.625,4200166.0,213
620842.4375,4206347.5,215
622382.4375,4208801.5,216
621438.6875,4207952.5,217
620432.1875,4207654.5,218
620705.6875,4210842.0,219
618233.1875,4211900.0,220
616444.4375,4210014.5,221
618958.625,4208111.5,222
615533.625,4208194.0,223
622302.4375,4213437.5,224
620175.875,4212240.5,225
618598.625,4212887.0,226
590536.0625,4213751.0,227
587980.5,4220547.5,228
588024.0,4221139.5,229
624352.0625,4211834.0,232
605623.9375,4235334.0,237
588033.4375,4215484.5,238
620171.75,4219633.5,239
615395.625,4219328.5,240
641895.8750000001,4208516.5,241
638683.1875,4211793.0,242
635133.625,4212840.0,243
633273.9375,4211326.5,244
631345.625,4214756.5,245
638817.875,4216453.0,246
635170.4375,4214520.5,247
634015.1875,4216437.5,248
632134.5625,4218603.5,249
632175.0,4217215.5,250
629827.75,4216585.5,251
627462.4375,4216463.5,252
631546.4375,4236310.5,253
631360.5,4235118.5,254
631571.5625,4233763.0,255
631426.1875,4233163.5,256
636535.8125,4235287.5,257
633314.3125,4235393.0,258
632552.375,4233660.0,259
631827.625,4232178.5,260
631905.5,4230359.0,261
633179.8125,4228466.5,262
632221.1875,4226976.5,263
631984.4375,4225284.5,264
631091.25,4223485.0,265
631070.0625,4222295.5,266
631289.5,4221229.0,267
631697.625,4219816.0,268
629256.8125,4220378.0,269
626871.1875,4219755.5,270
625126.625,4221403.5,271
624381.0,4219077.0,272
605245.75,4236976.5,273
637345.75,4229647.0,274
635542.125,4229615.0,275
636119.6875,4226160.0,276
634454.5625,4225637.5,277
637657.1875,4223313.5,278
634586.9375,4222445.5,279
630760.1875,4231768.0,280
630896.8125,4230314.5,281
630391.625,4229417.5,282
629403.0625,4229223.0,283
628928.625,4226857.5,284
628788.4375,4225515.5,285
627541.0625,4223149.5,286
626270.5,4222389.0,287
628872.0,4231936.0,288
627830.625,4231621.0,289
628130.4375,4230212.5,290
626822.375,4228235.0,291
624931.25,4226952.5,292
624074.0625,4224938.5,293
623763.125,4223037.0,294
623193.375,4221824.5,295
628905.5625,4252743.0,296
627633.3125,4250326.0,297
626433.9375,4247904.0,298
624725.5,4246059.0,299
623765.75,4243605.0,300
622700.5,4241281.0,301
621945.75,4238439.5,302
623262.8125,4237344.0,303
622416.0,4234913.0,304
622308.5,4232221.5,305
620526.0,4228156.0,306
618431.4375,4238744.5,307
618934.375,4236519.5,308
628051.0625,4269071.0,309
623344.9375,4266572.0,310
623488.0625,4259165.0,311
621997.6875,4254776.0,312
619911.4375,4248766.5,313
618262.25,4244148.5,314
616992.75,4236793.5,315
615935.375,4232392.0,316
616473.3125,4243967.0,317
616745.9375,4238622.5,318
614189.375,4243223.0,319
611470.875,4238825.0,320
614362.8125,4235236.5,321
614750.0625,4233770.0,322
615156.125,4233060.5,323
607124.0625,4235475.0,324
609429.0625,4235459.0,325
611764.3125,4234500.0,326
587823.0625,4224132.5,327
595501.8125,4215164.0,328
586524.5,4214278.5,329
629891.625,4272969.5,330
629038.9375,4269161.0,331
628650.75,4264609.5,332
626013.625,4261384.5,333
628614.125,4259463.5,334
628752.3125,4255115.0,335
629596.6875,4251881.0,336
629229.5,4249282.0,337
628130.5625,4245779.0,338
624538.25,4243096.5,339
624757.875,4240625.5,340
627726.25,4237278.5,341
630298.0,4234283.0,342
629777.75,4233513.5,343
626301.25,4233288.5,344
626242.8125,4229084.5,346
624212.8125,4227501.0,347
622026.3125,4224923.5,348
619570.375,4225750.5,349
616949.8125,4226701.0,350
614843.9375,4222528.5,351
613332.125,4218718.5,352
610418.25,4216250.5,353
605187.8125,4212988.5,354
601451.1875,4214097.0,355
597549.5,4211557.0,356
592570.8125,4212285.0,357
584737.8125,4213362.5,358
581339.1875,4212608.5,359
577182.6875,4210734.0,360
575688.9375,4209950.5,361
588514.0,4212713.0,362
585650.125,4216982.0,363
582403.25,4220726.0,364
582893.875,4218073.5,365
584113.9375,4215092.0,366
579898.5,4214940.0,367
584038.4375,4233013.5,368
575244.1875,4230363.0,369
575783.6875,4230210.0,370
584825.5625,4230665.5,371
584477.9375,4229699.5,372
584202.875,4227650.0,373
583405.8125,4226001.0,374
582029.375,4225318.5,375
582619.125,4223721.5,376
580409.6875,4221311.0,377
580883.9375,4219731.0,378
576604.75,4229434.5,379
577759.125,4227817.0,380
577905.1875,4224699.5,381
578714.3125,4223766.5,382
577161.8125,4227841.0,383
579006.0625,4218597.5,384
578711.375,4215837.5,385
579664.4375,4223945.0,386
581618.25,4227654.0,387
581275.0625,4226199.0,388
578504.25,4227633.0,389
580296.875,4226578.0,390
578493.0,4224914.5,391
582979.9375,4231027.0,392
581325.75,4228890.0,393
582795.625,4228606.0,394
586195.9375,4231292.5,395
577863.625,4230035.0,396
585056.9375,4228978.0,397
585043.4375,4227579.0,398
586624.5625,4226536.0,399
582672.125,4229113.0,400
593844.3125,4230098.5,403
588520.0,4231198.5,404
587355.0,4231297.5,405
594670.3125,4226141.0,406
596422.625,4231057.5,408
594540.0,4228496.5,409
595508.0625,4226568.5,410
595793.625,4225392.0,412
591665.6875,4226779.5,413
613242.9375,4216670.0,414
611898.25,4215672.5,416
597984.1875,4214857.0,417
597598.9375,4216803.5,418
595611.0,4221949.5,420
593356.0625,4224968.5,421
591322.6875,4225405.0,422
588523.875,4226635.5,425
583038.25,4223480.0,428
596047.125,4215896.5,432
593818.75,4216586.0,433
590875.5625,4218175.5,434
588576.0625,4218088.0,436
579851.875,4218954.0,440
578840.8125,4220274.0,442
579941.3125,4223084.5,443
579236.25,4219359.5,444
581392.125,4223626.5,445
637184.375,4235591.0,446
637278.9375,4235248.5,447
636405.4375,4238134.0,448
634454.1875,4236905.5,449
631203.1875,4242527.0,451
630151.0625,4241166.0,452
630697.6875,4239034.0,453
631451.125,4236935.0,454
630645.4375,4235900.5,455
650013.9375,4202023.5,456
648109.3750000001,4201934.0,457
606246.375,4211305.5,459
606661.5,4210815.5,460
608516.625,4209693.5,461
602421.1875,4211087.0,462
600739.9375,4209909.0,463
600535.5,4213950.5,464
599135.5,4212739.0,465
599892.6875,4211891.5,466
606637.5625,4209337.0,467
614667.625,4212004.0,469
604622.625,4211415.0,470
602828.625,4211026.0,471
639151.9171346205,4185391.2771015544,570
627310.8125,4273644.5,700
625291.125,4274900.0,701
624907.4375,4277948.5,702
622378.0625,4278190.5,703
623106.5,4259446.5,710
621738.8125,4255100.5,711
620010.875,4250018.0,712
618586.0625,4245934.0,713
617443.125,4240806.5,714
644784.282121603,4184263.4351714365,800
644293.6150041994,4184593.3093483397,801
643942.1912579511,4184822.0663152374,802
643158.4667838719,4185422.8523614863,803
642814.6472868258,4185436.8858103454,804
644439.9908879494,4183693.519852071,805
644077.4675266441,4184065.9966735775,806
643773.9230537417,4184636.5689910636,807
643102.9300083783,4185045.0987703833,808
642817.6438496355,4185124.978894831,809
642336.0808136774,4185252.787093948,810
640950.7312268219,4185218.552754899,811
640234.0923960598,4185026.8404562236,812
639147.6667574431,4183090.927823613,813
638620.422077507,4184427.0852266056,814
631626.3364237034,4183226.675730902,815
