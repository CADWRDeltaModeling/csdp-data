425
652083 4172133 1
652497.6 4174602 2
651897.1 4175821 3
650043.9 4176492 4
649492.2 4179509 5
649711.7 4182405 6
648587 4183898 7
647325.1 4185605 8
648462 4187495 9
647568.9 4189903 10
647605.5 4191853 11
647038.6 4195084 12
647812.8 4198071 13
647029.4 4198986 14
646377.2 4199992 15
645417.1 4200449 16
645889.5 4200936 17
646297.9 4201455 18
645194.5 4201851 19
644234.4 4202278 20
643310.9 4203131 21
642091.7 4204472 22
640567.7 4205569 23
639604.5 4206057 24
637614.2 4205996 25
636727.2 4206423 26
636861.3 4207764 27
635175.8 4207185 28
635468.4 4208221 29
634224.8 4209684 30
632496.6 4209959 31
632719.1 4210782 32
630125.2 4212549 34
628704.9 4212763 35
628756.7 4214104 36
625717.8 4214835 38
625224.1 4215902 39
625013.7 4216938 40
621572.5 4217883 41
618984.8 4216237 42
615717.3 4215719 43
615796.6 4213128 44
611690.9 4209745 45
607033.6 4208313 46
602723.7 4209471 47
646611.9 4186215 48
646166.9 4187099 49
645462.8 4187068 50
644411.2 4186733 51
643115.8 4187038 52
642695.2 4186794 53
641753.4 4185666 54
639287.5 4185818 56
639147.3 4184965 57
639183.9 4184477 58
637909.8 4184233 59
637157 4184721 60
635815.9 4184752 61
634916.7 4184264 62
634255.3 4183258 63
633505.5 4182496 64
632444.8 4182405 65
631496.8 4183258 66
629951.5 4184203 67
629216.9 4184934 68
628357.4 4185514 69
627025.4 4186215 70
627571 4187160 71
627482.6 4187617 72
627141.2 4188592 73
626854.7 4189476 74
626525.5 4190512 75
626004.3 4191061 76
625586.8 4191640 77
625199.7 4192829 78
625333.8 4194078 79
626095.8 4194810 80
625583.7 4195846 81
626388.4 4196883 82
626178.1 4197218 83
627095.5 4197888 84
626918.7 4198925 85
626565.2 4199900 86
626815.1 4200601 87
625876.3 4200357 88
626318.3 4201424 89
625272.8 4201546 90
626172 4202034 91
625489.2 4202552 92
625147.9 4203558 93
624675.4 4204564 94
624742.5 4205295 95
625227.1 4205844 96
624812.6 4206240 97
624772.9 4207246 99
626754.1 4208496 100
624657.1 4210050 102
624498.6 4213342 103
642091.7 4187830 104
642670.8 4189964 105
642914.6 4191335 106
642274.6 4193134 107
641134.6 4194200 108
639388.1 4194383 109
637955.5 4194810 110
636748.5 4194048 111
634785.6 4193652 112
632947.7 4194322 113
632353.3 4195328 114
632069.9 4196029 115
631198.1 4196334 116
630561.1 4197157 117
630228.9 4197736 118
629399.8 4198071 119
629469.9 4199108 120
628973.1 4199870 121
628829.8 4200784 122
629704.6 4200845 123
629177.3 4201973 124
628814.6 4203192 125
628802.4 4204167 126
628823.7 4205112 127
629207.8 4205996 128
629951.5 4206789 129
630750.1 4206880 130
630966.5 4207673 131
630283.7 4207734 132
630235 4208983 133
629259.6 4211361 134
630491 4204320 135
627150.4 4213007 37
643103.6 4200693 138
642442.2 4202186 139
635584.2 4205630 140
634127.3 4204807 141
634041.9 4203497 142
632493.5 4203466 143
631207.3 4203466 144
629890.5 4203436 145
637906.8 4199534 146
636017 4201638 147
634584.5 4202613 148
643076.2 4181064 154
642305 4181338 155
642027.7 4182069 156
641469.9 4181643 157
640104.4 4182222 159
639644.1 4182862 160
639382 4183471 149
648961.9 4180271 162
646925.8 4181947 163
645450.6 4183624 164
643597.4 4184843 165
645411 4183014 166
643597.4 4184508 167
641622.3 4185209 168
639635 4184965 169
640415.3 4186794 170
638324.4 4186763 171
636541.3 4186702 172
635770.1 4186672 173
634453.4 4186641 174
633423.2 4186641 175
632246.6 4186611 176
630990.9 4186580 177
628921.3 4186550 178
625556.3 4186093 179
625181.4 4185636 180
624666.3 4184020 181
628439.7 4188318 182
628845.1 4189354 183
629037.1 4189903 184
628418.4 4189964 185
628454.9 4190756 186
627787.4 4190482 187
632021.1 4193804 188
630619 4193012 189
629759.5 4192554 190
628933.5 4192097 191
627400.3 4191183 192
623861.6 4187922 193
629073.7 4196974 194
627589.3 4196944 195
625218 4197462 196
624117.6 4197675 197
622618 4197340 198
622422.9 4198559 199
622230.9 4199717 200
622401.6 4201363 201
622782.6 4202491 202
623569 4203375 203
622654.6 4203893 204
621066.6 4204015 205
619463.3 4203802 206
628765.8 4207154 207
627129.1 4207703 208
623041.7 4188562 209
623965.2 4188958 210
624559.6 4189750 211
625019.8 4191091 212
627586.3 4199900 213
621066.6 4204320 214
620981.2 4206118 215
622377.2 4208435 216
621542.1 4207703 217
620481.4 4207429 218
621380.5 4210020 219
618308.1 4211665 220
616528.1 4209806 221
619054.9 4207916 222
615546.7 4208130 223
622621.1 4213220 224
620274.1 4212001 225
618683 4212610 226
590632.3 4213555 227
621270.8 4212580 230
623950 4212885 231
624251.7 4211513 232
621395.8 4210782 234
622520.5 4211513 235
615613.7 4207977 236
612416.4 4208191 237
588166.5 4215232 238
620268 4219438 239
615491.8 4219133 240
641975.9 4208282 241
638732.8 4211604 242
635255 4212580 243
633481.1 4211239 244
631442 4214561 245
638958.3 4216298 246
635273.3 4214287 247
634206.5 4215994 248
632313.7 4218310 249
632219.2 4216847 250
629924.1 4216390 251
627558.8 4216268 252
631646.2 4236019 253
631448.1 4234891 254
631634 4233520 255
631481.6 4232819 256
636648 4235074 257
633423.2 4235196 258
632688.6 4233428 259
632005.9 4231904 260
631987.6 4230106 261
633276.9 4228216 262
632365.5 4226753 263
632143 4224955 264
631201.2 4223278 265
631112.8 4222090 266
631393.2 4220962 267
631795.5 4219529 268
629363.2 4220139 269
626967.5 4219560 270
624913.2 4220962 271
624443.8 4218828 272
605341.9 4236781 273
635660.4 4229374 275
634550.9 4225442 277
637605 4223034 278
634630.2 4222212 279
630856.8 4231538 280
631024.4 4230106 281
630487.9 4229222 282
629241.3 4228551 283
629024.9 4226662 284
628884.7 4225320 285
627665.5 4222913 286
626336.6 4222181 287
629015.8 4231660 288
627936.8 4231356 289
628269 4230014 290
626949.2 4228033 291
625065.6 4226692 292
624178.6 4224741 293
623876.8 4222821 294
623255 4221602 295
628835.9 4252448 296
627729.5 4250131 297
626516.4 4247693 298
624821.7 4245864 299
623849.4 4243365 300
622816.1 4241048 301
622041.9 4238244 302
623364.8 4237147 303
622517.4 4234678 304
622404.7 4232026 305
620719.1 4227942 306
628147.1 4268876 309
623441 4266377 310
623584.2 4258970 311
622093.8 4254581 312
619810.8 4248607 313
617088.9 4236598 315
616113.6 4231965 316
616579.9 4243700 317
616842.1 4238427 318
614278.7 4242938 319
611678.7 4238427 320
614421.9 4235013 321
614827.3 4233520 322
615363.8 4232880 323
607225.6 4235196 324
609231.2 4235105 325
611526.3 4235013 326
587840.3 4223796 327
594195.4 4214073 328
586794.9 4213982 329
630000.3 4272686 330
629006.6 4268968 331
628720.1 4264396 332
625730 4261957 333
628628.7 4259214 334
630719.6 4255526 335
628479.3 4253697 336
629284 4249034 337
628360.4 4245742 338
624623.6 4242877 339
624840 4240378 340
627778.3 4237055 341
630402.6 4234038 342
629860.1 4233245 343
626397.5 4233093 344
626370.1 4230807 345
626367.1 4228917 346
624163.3 4227119 347
622139.5 4224680 348
619682.8 4225503 349
616832.9 4226082 350
614940.1 4222333 351
613428.3 4218523 352
610514.4 4216055 353
605284 4212793 354
601172.3 4213860 355
597645.7 4211361 356
592397.1 4212519 357
585740.3 4212946 358
581119.5 4212184 359
577279 4210538 360
575950.1 4209532 361
588596.2 4212366 362
585746.4 4216786 363
582841.6 4220261 364
582728.8 4218676 365
584210.2 4214896 366
579994.8 4214744 367
584798.4 4218645 368
575340.5 4230167 369
575880 4230014 370
584947.8 4230411 371
584454 4229557 372
584301.6 4227332 373
583414.6 4225839 374
582152.8 4225046 375
582649.6 4223522 376
580485.5 4221053 377
581192.6 4219499 378
576623.7 4229252 379
577867.3 4227606 380
577916 4224498 381
578784.7 4223522 382
579333.4 4221267 383
579077.3 4218402 384
578821.3 4215628 385
579827.1 4223705 386
581527.9 4227149 387
581381.6 4225961 388
579034.7 4226631 389
580418.5 4226387 390
578510.4 4224711 391
583192.1 4231264 392
581454.8 4228612 393
582884.3 4228368 394
586276.7 4231081 395
578236.1 4230868 396
585142.9 4228734 397
585136.8 4227332 398
586767.4 4226326 399
586490.1 4226052 401
584685.7 4226022 402
593951.6 4229892 403
588642 4230959 404
587453.2 4231081 405
594817.2 4225930 406
596514.9 4230898 408
594872.1 4228308 409
595655.4 4226265 410
595792.6 4225229 412
591769.2 4226509 413
598014.6 4215384 415
598072.5 4214652 417
597843.9 4216237 418
595707.2 4221754 420
593451.7 4224650 421
591397.3 4225138 422
588614.5 4226479 425
583183 4223187 428
593915 4216390 433
591613.8 4216725 434
588666.3 4217822 436
579888.1 4219956 438
579879 4218737 440
578937.1 4220078 442
580022.2 4222821 443
579318.1 4219164 444
581460.9 4223339 445
637227.1 4235287 446
637345.9 4235013 447
636501.7 4237939 448
634538.7 4236659 449
630984.8 4242877 450
631295.7 4242267 451
630262.4 4240804 452
630795.8 4238793 453
631566.9 4236720 454
630759.2 4235623 455
625742.2 4206636 98
630658.6 4205265 136
631253 4205935 137
619030.5 4236324 308
618527.6 4238549 307
631593.8 4211665 33
625072.9 4211397 101
618358.4 4243953 314
