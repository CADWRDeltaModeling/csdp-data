;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      427
586698.625,4214178.0,329
594099.1875,4214269.0,328
587744.0,4223991.5,327
611430.1875,4235208.5,326
609135.125,4235300.5,325
607129.5,4235391.5,324
615267.6875,4233075.5,323
614731.1875,4233715.5,322
627840.5625,4231551.5,289
614325.8125,4235208.5,321
628919.5625,4231855.5,288
611582.625,4238622.5,320
626240.3125,4222376.5,287
627569.1875,4223108.5,286
628788.4375,4225515.5,285
628928.625,4226857.5,284
629145.0,4228746.5,283
630391.625,4229417.5,282
630928.125,4230301.5,281
630760.5625,4231733.5,280
614182.5625,4243133.5,319
616745.9375,4238622.5,318
616483.75,4243895.5,317
616017.4375,4232160.5,316
616992.75,4236793.5,315
618262.25,4244148.5,314
619714.6875,4248802.0,313
621997.6875,4254776.0,312
634533.875,4222407.5,279
623488.0625,4259165.0,311
637508.625,4223229.5,278
623344.9375,4266572.0,310
634454.5625,4225637.5,277
635564.125,4229569.5,275
605245.75,4236976.5,273
624347.5,4219023.5,272
624816.9375,4221157.5,271
626871.1875,4219755.5,270
628051.0625,4269071.0,309
618934.375,4236519.5,308
618431.4375,4238744.5,307
620622.875,4228137.5,306
622308.5,4232221.5,305
622421.1875,4234873.5,304
623268.625,4237342.5,303
621945.75,4238439.5,302
629266.875,4220334.5,269
622719.9375,4241243.5,301
631699.125,4219724.5,268
623753.25,4243560.0,300
631296.875,4221157.5,267
631016.4375,4222285.5,266
631104.875,4223473.5,265
632046.6875,4225150.5,264
632269.1875,4226948.5,263
633180.625,4228411.5,262
631891.3125,4230301.5,261
631909.625,4232099.5,260
632592.3125,4233623.5,259
633326.9375,4235391.0,258
636551.75,4235269.0,257
631385.3125,4233014.5,256
631537.75,4233715.5,255
631351.875,4235086.5,254
631549.9375,4236214.0,253
627462.4375,4216463.5,252
629827.75,4216585.5,251
632122.8125,4217042.5,250
632217.3125,4218505.5,249
634110.125,4216189.5,248
635176.875,4214482.5,247
638861.875,4216493.5,246
631345.625,4214756.5,245
633384.6875,4211434.5,244
635158.5625,4212775.5,243
638636.375,4211799.5,242
641879.4375,4208477.5,241
615395.625,4219328.5,240
620171.75,4219633.5,239
588070.25,4215428.0,238
612320.1875,4208386.5,237
615517.5,4208172.5,236
622424.1875,4211708.5,235
621299.5,4210977.5,234
624155.375,4211708.5,232
622326.5625,4198754.5,199
623853.6875,4213080.5,231
622521.6875,4197535.5,198
621174.5,4212775.5,230
624021.25,4197870.5,197
625121.625,4197657.5,196
627492.9375,4197139.5,195
628977.3125,4197169.5,194
623765.25,4188117.75,193
627303.9375,4191378.75,192
628837.125,4192292.75,191
629663.125,4192749.75,190
587707.8979938272,4220110.2968107,228
590536.0625,4213751.0,227
618586.75,4212805.5,226
620177.8125,4212196.5,225
622524.8125,4213415.5,224
615450.5,4208325.5,223
618958.625,4208111.5,222
630522.625,4193207.75,189
616431.875,4210001.5,221
631924.6875,4193999.5,188
618211.875,4211860.5,220
627691.0,4190677.75,187
628358.5,4190951.75,186
628322.0,4190159.75,185
628940.75,4190098.75,184
628748.75,4189549.7500000005,183
628343.3125,4188513.75,182
624569.9375,4184215.7500000005,181
625085.0625,4185831.75,180
621284.1875,4210215.5,219
620385.125,4207624.5,218
621445.8125,4207898.5,217
622280.875,4208630.5,216
620884.875,4206313.5,215
620970.3125,4204515.5,214
627489.9375,4200095.5,213
624923.4375,4191286.75,212
625459.9375,4186288.75,179
624463.25,4189945.75,211
628824.9375,4186745.75,178
623868.875,4189153.75,210
630894.5,4186775.7499999995,177
632150.1875,4186806.75,176
633326.8125,4186836.75,175
634357.0,4186836.5,174
635673.6875,4186867.4999999995,173
636554.0,4186941.0,172
638228.0,4186958.5,171
640318.8749999999,4186989.5,170
622945.375,4188757.75,209
627032.6875,4207898.5,208
628669.375,4207349.5,207
619367.0,4203997.5,206
620970.3125,4204210.5,205
622558.25,4204088.5,204
623472.6875,4203570.5,203
622686.25,4202686.5,202
639538.6249999999,4185160.5,169
622305.25,4201558.5,201
641525.875,4185404.5,168
622134.5625,4199912.5,200
643501.0,4184703.5,167
645314.6250000001,4183209.5,166
643501.0,4185038.5,165
645354.1875,4183819.4999999995,164
646829.375,4182142.5000000005,163
648865.5,4180466.5,162
639547.6875,4183057.4999999995,160
640008.0,4182417.5,159
641373.5,4181838.5,157
641931.3125,4182264.5,156
642208.625,4181533.4999999995,155
642979.8125,4181259.5000000005,154
639285.625,4183666.5000000005,149
634488.0625,4202808.5,148
635920.5625,4201833.5,147
637810.375,4199729.5,146
629794.0625,4203631.5,145
631110.875,4203661.5,144
632397.0625,4203661.5,143
633945.4375,4203692.5,142
634030.875,4205002.5,141
635487.75,4205825.5,140
642345.75,4202381.5,139
643007.125,4200888.5,138
631156.5625,4206130.5,137
630562.1875,4205460.5,136
630394.5625,4204515.5,135
629163.1875,4211556.5,134
630138.5625,4209178.5,133
630187.25,4207929.5,132
630870.0625,4207868.5,131
630653.6875,4207075.5,130
629855.0625,4206984.5,129
629111.375,4206191.5,128
628727.3125,4205307.5,127
628706.0,4204362.5,126
628718.1875,4203387.5,125
629080.875,4202168.5,124
629608.1875,4201040.5,123
628733.375,4200979.5,122
628876.6875,4200065.5,121
629373.5,4199303.5,120
629303.375,4198266.5,119
630132.5,4197931.5,118
630464.6875,4197352.5,117
631101.6875,4196529.5,116
631973.5,4196224.5,115
632256.875,4195523.5,114
632851.3125,4194517.5,113
634689.1875,4193847.5,112
636652.0625,4194243.4999999995,111
637859.0625,4195005.5,110
639291.6875,4194578.5,109
641038.1875,4194395.5,108
642178.1875,4193329.5,107
642818.1875,4191530.5,106
642574.375,4190159.5000000005,105
641995.3124999999,4188025.5,104
624402.3125,4213537.5,103
624560.75,4210245.5,102
624976.5625,4211592.5,101
626657.75,4208691.5,100
624676.5625,4207441.5,99
625645.8125,4206831.5,98
624716.25,4206435.5,97
625130.75,4206039.5,96
624646.125,4205490.5,95
624579.0625,4204759.5,94
625051.5625,4203753.5,93
625392.8125,4202747.5,92
626075.625,4202229.5,91
625176.4375,4201741.5,90
630662.9375,4235818.5,455
631470.6875,4236915.0,454
630699.5625,4238988.0,453
630166.1875,4240999.0,452
631199.5,4242462.0,451
630888.5625,4243072.0,450
626221.9375,4201619.5,89
625779.9375,4200552.5,88
626718.75,4200796.5,87
626468.8125,4200095.5,86
626822.3125,4199120.5,85
626999.125,4198083.5,84
626081.75,4197413.5,83
626292.0,4197078.5,82
634442.4375,4236854.0,449
625487.3125,4196041.5,81
636405.4375,4238134.0,448
625999.4375,4195005.5,80
637249.625,4235208.0,447
637130.8125,4235482.0,446
581364.625,4223535.0,445
579221.8125,4219360.0,444
579925.875,4223017.0,443
578840.8125,4220274.0,442
579782.6875,4218933.0,440
625237.4375,4194273.75,79
625103.3125,4193024.75,78
625490.4375,4191835.7500000005,77
625907.9375,4191256.75,76
626429.125,4190707.75,75
626758.3125,4189671.75,74
627044.8125,4188787.7500000005,73
627302.0,4187963.0,72
627474.625,4187355.75,71
579791.8125,4220152.0,438
626929.0625,4186410.7499999995,70
588570.0,4218018.0,436
591517.5625,4216921.0,434
593818.75,4216586.0,433
586671.125,4226521.5,399
585040.5,4227527.5,398
585046.625,4228929.5,397
578508.9869422007,4227748.015545141,396
586180.4375,4231276.5,395
582788.0,4228564.0,394
581358.5,4228808.0,393
583095.8125,4231460.0,392
578414.125,4224907.0,391
580322.1875,4226583.0,390
628267.0,4185764.0,69
629120.5,4185129.75,68
629855.125,4184398.75,67
631400.4375,4183453.7500000005,66
632348.4375,4182600.7499999995,65
633409.125,4182691.7500000005,64
634158.9375,4183453.7500000005,63
634820.3125,4184459.75,62
635719.5,4184947.5,61
583086.6875,4223383.0,428
637060.625,4184916.5,60
588518.25,4226674.5,425
591301.0625,4225333.5,422
578938.375,4226827.0,389
593355.4375,4224845.5,421
581285.3125,4226157.0,388
595611.0,4221949.5,420
581431.625,4227345.0,387
579730.8125,4223901.0,386
578725.0,4215824.0,385
578981.0,4218598.0,384
579237.125,4221463.0,383
578688.375,4223718.0,382
577819.6875,4224694.0,381
577771.0,4227802.0,380
637813.4375,4184428.5000000005,59
639087.5,4184672.5,58
639050.875,4185160.5,57
639191.125,4186013.5,56
641657.0,4185861.4999999995,54
642598.8125,4186989.5,53
643019.375,4187233.5,52
644314.8125,4186928.5,51
597598.9375,4216803.5,418
645366.375,4187263.5,50
597976.3125,4214847.5,417
597918.375,4215579.5,415
591672.9375,4226704.5,413
595696.375,4225424.5,412
576527.375,4229448.0,379
581096.3125,4219695.0,378
595559.1875,4226460.5,410
580389.1875,4221249.0,377
582553.3125,4223718.0,376
582056.5,4225242.0,375
583318.3125,4226035.0,374
584205.3125,4227528.0,373
584357.6875,4229752.5,372
584851.5,4230606.5,371
575783.6875,4230210.0,370
646070.5,4187294.5,49
646515.5000000001,4186410.5,48
602627.5,4209666.5,47
606937.4375,4208508.5,46
611594.75,4209940.5,45
615700.375,4213323.5,44
615621.125,4215914.5,43
618888.5625,4216432.5,42
594775.875,4228503.5,409
621476.25,4218078.5,41
596418.6875,4231093.5,408
624917.375,4217133.5,40
594721.0,4226125.5,406
587356.9375,4231276.5,405
588545.75,4231154.5,404
593855.375,4230087.5,403
584589.4375,4226218.0,402
575244.1875,4230363.0,369
586393.8125,4226247.5,401
583961.4892489712,4233078.634773662,368
582655.75,4229097.5,400
579898.5,4214940.0,367
584113.9375,4215092.0,366
582632.5,4218872.0,365
582745.3125,4220457.0,364
585650.125,4216982.0,363
588499.9375,4212562.0,362
575853.8125,4209728.0,361
577182.6875,4210734.0,360
625127.8125,4216097.5,39
625621.5,4215030.5,38
627054.0625,4213202.5,37
628660.3125,4214299.5,36
628608.5,4212958.5,35
630028.8125,4212744.5,34
631497.375,4211860.5,33
632622.6875,4210977.5,32
632400.1875,4210154.5,31
634128.375,4209879.5,30
581023.1875,4212380.0,359
585644.0,4213142.0,358
592300.875,4212715.0,357
597549.5,4211557.0,356
601076.125,4214055.5,355
605187.8125,4212988.5,354
610418.25,4216250.5,353
613332.125,4218718.5,352
614843.9375,4222528.5,351
616736.75,4226277.5,350
635371.9375,4208416.5,29
635079.3125,4207380.5,28
636764.8125,4207959.5,27
636630.75,4206618.5,26
637517.75,4206191.5,25
639508.0,4206252.5,24
640471.25,4205764.5,23
641995.25,4204667.5,22
643214.4374999999,4203326.5,21
644137.9375,4202473.5,20
619586.625,4225698.5,349
648365.5625,4187690.5,9
622043.25,4224875.5,348
624067.0625,4227314.5,347
647151.0,4185852.0,8
648490.5624999999,4184093.5,7
626270.875,4229112.5,346
649615.3124999999,4182600.5,6
626273.875,4231002.5,345
649395.8125,4179704.5,5
626301.25,4233288.5,344
649947.5,4176687.5000000005,4
629763.875,4233440.5,343
651800.6875,4176016.25,3
630298.0,4234283.0,342
652401.1875000001,4174797.25,2
627682.0625,4237250.5,341
651986.625,4172328.2500000005,1
624743.8125,4240573.5,340
645098.0,4202046.5,19
646201.4374999999,4201650.5,18
645793.0,4201131.5,17
645320.625,4200644.5,16
646280.75,4200187.5,15
646932.9375,4199181.5,14
647716.3125,4198266.5,13
646942.125,4195279.5,12
647509.0625,4192048.5000000005,11
647472.4375,4190098.5,10
624527.4375,4243072.0,339
628264.1875,4245937.0,338
629187.8125,4249229.0,337
628383.125,4253892.0,336
630623.4375,4255721.0,335
628532.5625,4259409.0,334
625633.875,4262152.0,333
628624.0,4264591.0,332
624725.5,4246059.0,299
628910.5625,4269163.0,331
626420.25,4247888.0,298
629904.25,4272881.0,330
627633.3125,4250326.0,297
628739.75,4252643.0,296
623158.75,4221797.5,295
623780.5625,4223016.5,294
624082.375,4224936.5,293
624969.375,4226887.5,292
626852.9375,4228228.5,291
628172.75,4230209.5,290
