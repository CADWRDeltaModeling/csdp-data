;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      22
615374.3299287185,4219538.540395569,7_mile@3_mile
621519.3229452168,4218672.1768282885,7_mile@sjr
616015.4920929506,4213273.557979698,FalseBarrier
627294.7192011583,4187980.382940997,clifton_court
613242.4440624218,4216675.39407366,decker_is_north_weir
611895.640197218,4215686.524569028,decker_is_south_weir
630345.27712,4234274.740411251,delta_cross_channel
578827.3915500746,4215030.450602861,goodyear_sl
636502.2348807644,4186975.304674783,grant_line_barrier
634765.9481673968,4193868.910057635,middle_r_barrier
597590.1092166901,4216811.2200855035,montezuma_salinity_control
581715.7265187072,4218892.239519224,morrow_c_line_outfall
580739.4462395692,4219610.781804669,morrow_m_line_outfall
579267.2155786289,4218747.75003791,morrow_sys_intake
647196.1886412773,4185854.2862227494,old_r@head_barrier
628262.7615905908,4185770.630953449,old_r@tracy_barrier
649386.6688098945,4179709.5160144614,paradise_cut_weir
597540.7275429484,4216707.080714259,roaring_river_slough_intake
620974.3523706995,4204346.447983768,sandmound_sl
639260.5287332154,4183738.337926453,tom_paine_sl
588121.643232379,4220599.255807898,tule_red_weirs
618569.0787308341,4245952.57608175,yolo_flyway_weir
