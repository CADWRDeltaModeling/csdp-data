﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      149
576633.3,4211159,BENBR
600859.1,4214643.6,CSE
579121.895,4214883,FLT
624614.6,4207543.5,HLL
630737.3,4207200.2,HLT2
616731,4217465,TWI
640088,4185530,OTWW
635798.2,4185059.9,TWA
612410.9,4210203.7,BLP
610748.9,4216702.8,SDI
629219.1,4233351.8,GES
615180.4,4216618.4,SR3
629664.2,4235427.1,SDC
605228,4237166.9,BKS
612908.6,4237177.1,UCS
615105,4224350,RVB
627243.2,4188117.2,WCI
628839.5,4200455,MDM
615252.9,4224292.9,RIV
624476.9,4208582.2,HOL2
616657.3,4235072.2,DWS
632927.2,4194823.6,VIC
627753,4186838.8,GLC2
617644.9,4226137.5,SOI
630645,4183522,WCNM
623124,4259467.4,LIS
643018.6,4187320.1,UNI
629247.7,4247651,CCW
580303.5,4226742.3,SNC
615115,4233613,LIB
649512,4179437,DVI
628839.5,4200455,MDMZQ
625540.70,4217496.70,SAL
597238.3,4211183.7,PTS
582994.8199,4223547.67,HUN
627898.6,4185906.3,OBD
620996.1,4210486.7,BET2
643589.2414,4184870.011,PCSB
577650.9,4223639,IBS
580533.214,4219949.694,GOD
625274.8,4218552.5,MOK2
615196.3,4218095.3,TSL
615192.5278,4218085.215,TSS
619885.2,4204031,RSL
594757.5,4211123.3,MAL
597451.6,4219938,NSL
629804,4184307,MHCM
628312.5,4185763.1,OAD
623525.5,4259677.4,CM72
613995.8,4206152.6,CNT
621194.1,4204133.5,RSD
584309.0232,4220037.891,GZL
608116.21,4215165.61,M13
591743.04,4212444.61,C24
653005.8,4171637.9,VER
605075.1,4208474.7,ANC
643575.2,4202944.9,RRI
635762.3,4206110.6,TRN
586986.9,4219943,GZB
610598.8,4215917.6,EMM
619281.8,4227913.6,SXS
626573,4213393.1,PRI
620970,4251599.2,CM66
636491.6,4185281.5,OLD
633766.8116,4183139.204,ORFU
618511,4244595,CM62
579253,4219416,GYS
638631.8,4186457.6,DGL
616676.6,4208098.2,DSJ
602123.11,4213753.24,CO5
618409.8,4245456.2,LBTOE
583902.55,4213517.57,C16
605282.66,4213133.12,C10
630172.109,4186906.468,GLW
580045,4225811,TEA
615024.3,4212414.2,JER
579678,4223160,CYG
600858.7,4214644.1,CLL
619475.5,4208005.7,FRP
639555,4185573,PCCU
637754.4,4187026.5,GLE
629874.3,4233686.1,SWE
630666.9,4231648.1,MKN
632231.1776,4182733.49,OAAD
623008.4,4211892.7,FRK
626952,4187911.6,CLC
629291.6,4192502.2,VCU
653005.8,4171637.9,SJR
645200.2,4181269.9,TPP
647576.1,4186166.1,SJL
639072,4185270,PCCD
597605.9,4211894.6,CONFL
643229,4184985,PDUP
646735.2,4199969.7,SJG
639228.5,4183752.9,TPI
627213.4,4213060.7,PPT
648060.2,4187435.7,SJD
583348,4226330,VOL
639778,4185041,PDC
585550.4,4212803.2,PCT
631868.1,4217577.6,LPS
567940.8,4212900.6,CARQB
631678,4183047,OBRD
647500.8,4192114.6,BDT
622318.4,4234477.5,SUS
639164.7,4183509.3,SUR
590134.7,4227040.1,BDL
630762.5,4257477,FPT
616742.9,4232844.4,MIR
643723.1587,4185003.321,PCNB
625994.6,4209807.9,ORQ2
631586.4,4219845,STI
618521.7,4214201.8,FCT
593045.1,4214379.2,HON
624652.3,4214658.4,OSJ2
642469,4181997,TPPA
642184.4,4193313.5,MHO
637086,4184987,OTBD
623598.2,4238356.2,SSS
625718.9,4194688.9,OH4
613974.4,4218374.1,TMS
614250.8,4241943.7,SGG
616952.5,4212848.6,FAL2
649126.1,4183436.8,MSD2
635780.8,4193802,MTB
638981.8,4184006.2,SGA
608608.2,4214765.6,SSI
617515.3,4228186.2,RYF
617515,4228186,RYE
582761,4218277.6,GRIZZB
588041.6,4215616.3,RYC
597578.3032,4216762.676,MSL
614797.6,4223035.8,SRV
625718.9,4194688.9,OH4
623426.6,4202761.2,WDCUT
639210.2727,4181357.384,DAR
647096.2,4185827.7,OH1
642021.8,4186071.2,ORX
629727.3,4233179.3,GSS
629247.7,4247651,SRH
575432.5,4209227.7,MRZ
625406.5,4203423.6,BAC
634779.4549,4193764.353,MRX
642052.7,4188617.1,MRU
626882.7,4186454,DMC
630537,4183977,ORM
627377.4,4187715.2,ORI
584692.1,4227881.3,FMB
624631.5,4203880,HOLM
