﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      2628862.03,4200697.37,MDM_FLOW_144
628978.37,4200707.22,MDM_FLOW_145
