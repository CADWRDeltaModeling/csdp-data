﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      28
619734.2,4239063.4,HWB
630802.2,4234030.6,DLC
624348.3,4243212.4,SUT
615196.3,4218095.3,TSL
624476.9,4208582.2,HOL
625718.9,4194688.9,OH4
647096.2,4185827.7,OH1
630762.5,4257477,FPT
616952.5,4212848.6,FAL
636454.1,4186988.1,GCT
616676.6,4208098.2,DSJ
623598.2,4238356.2,SSS
629291.6,4192502.2,VCU
625222.5,4203213.9,OBI
629664.2,4235427.1,SDC
615024.3,4212414.2,JER
628084.5,4186853.4,GLC
635762.3,4206110.6,TRN
643575.2,4202944.9,RRI
618521.7,4214201.8,FCT
629727.3,4233179.3,GSS
597451.6,4219938,NSL
647500.8,4192114.6,BDT
625274.8,4218552.5,MOK
630093.3,4208185,HLT
639778,4185041,PDC
614797.6,4223035.8,SRV
629219.1,4233351.8,GES
