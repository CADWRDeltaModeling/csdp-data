;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      30
647500.8,4192114.6,BDT
620980,4210523,BET
626952,4187911.6,CLC
600858.7,4214644.1,CLL
610598.8,4215917.6,EMM
624614.6,4207543.5,HLL
615024.3,4212414.2,JER
594757.5,4211123.3,MAL
636491.6,4185281.5,OLD
585550.4,4212803.2,PCT
643018.6,4187320.1,UNI
629291.6,4192502.2,VCU
626882.7,4186454,DMC
625406.5,4203423.6,BAC
605228,4237166.9,BKS
613974.4,4218374.1,TMS
630666.9,4231648.1,NMR
631586.4,4219845,STI
615105,4224350,RVB
629727.3,4233179.3,GSS
597451.6,4219938,NSL
590134.7,4227040.1,BDL
583348,4226330,VOL
580303.5,4226742.3,SNC
577650.9,4223639,IBS
579253,4219416,GYS
625718.9,4194688.9,OH4
619885.2,4204031,RSL
605075.1,4208474.7,ANH
625540.70,4217496.70,SAL
