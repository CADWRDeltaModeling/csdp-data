;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype: landmark
;NumElements: 426
651986.618,4172328.340,1
652401.212,4174797.348,2
651800.711,4176016.365,3
649947.514,4176687.399,4
649395.808,4179704.424,5
649615.294,4182600.416,6
648490.589,4184093.431,7
648365.574,4187690.427,9
647472.465,4190098.435,10
647509.056,4192048.431,11
646942.144,4195279.431,12
647716.329,4198266.416,13
646932.927,4199181.423,14
646280.725,4200187.428,15
645320.626,4200644.437,16
645793.022,4201131.431,17
646201.419,4201650.425,18
645098.021,4202046.436,19
644137.922,4202473.445,20
643214.422,4203326.452,21
641995.221,4204667.459,22
640471.222,4205764.470,23
639508.023,4206252.477,24
637517.730,4206191.496,25
636630.732,4206618.502,26
636764.838,4207959.489,27
635079.340,4207380.510,28
635371.946,4208416.497,29
634128.361,4209879.494,30
632400.170,4210154.507,31
632622.675,4210977.497,32
630028.810,4212744.499,34
628608.529,4212958.507,35
628660.337,4214299.493,36
625621.478,4215030.506,38
625127.790,4216097.498,39
624917.399,4217133.489,40
621476.243,4218078.502,41
618888.565,4216432.537,42
615621.102,4215914.565,43
615700.391,4213323.592,44
611594.732,4209940.659,45
606937.439,4208508.715,46
602627.517,4209666.745,47
646515.483,4186410.455,48
646070.481,4187294.460,49
645366.382,4187263.469,50
644314.786,4186928.485,51
643019.388,4187233.502,52
642598.790,4186989.509,53
641656.996,4185861.526,54
639191.101,4186013.560,56
639050.905,4185160.565,57
639087.506,4184672.567,58
637813.410,4184428.586,59
637060.610,4184916.595,60
635719.513,4184947.614,61
634820.316,4184459.630,62
634158.921,4183453.644,63
633409.125,4182691.659,64
632348.428,4182600.676,65
631400.427,4183453.680,66
629855.128,4184398.684,67
629120.528,4185129.684,68
626929.033,4186410.690,70
627474.630,4187355.682,71
627044.831,4188787.677,73
626758.331,4189671.675,74
626429.132,4190707.671,75
625907.935,4191256.672,76
625490.437,4191835.671,77
625103.340,4193024.668,78
625237.439,4194273.660,79
625999.433,4195005.652,80
625487.336,4196041.650,81
626292.029,4197078.639,82
626081.731,4197413.638,83
626999.122,4198083.629,84
626822.322,4199120.624,85
626468.825,4200095.621,86
626718.722,4200796.616,87
625779.932,4200552.624,88
626221.926,4201619.615,89
625176.438,4201741.622,90
626075.628,4202229.613,91
625392.835,4202747.615,92
625051.539,4203753.612,93
624579.045,4204759.610,94
624646.144,4205490.605,95
625130.738,4206039.599,96
624716.243,4206435.600,97
624676.548,4207441.591,99
626657.728,4208691.564,100
624560.765,4210245.563,102
624402.285,4213537.530,103
641995.287,4188025.514,104
642574.377,4190159.499,105
642818.171,4191530.492,106
642178.165,4193329.494,107
641038.164,4194395.505,108
639291.668,4194578.525,109
637859.070,4195005.541,110
636652.077,4194243.559,111
634689.183,4193847.585,112
632851.286,4194517.604,113
632256.884,4195523.605,114
631973.483,4196224.604,115
631101.688,4196529.610,116
630464.691,4197352.609,117
630132.493,4197931.608,118
629303.400,4198266.612,119
629373.497,4199303.606,120
628876.700,4200065.605,121
628733.400,4200979.601,122
629608.190,4201040.594,123
629080.894,4202168.592,124
628718.195,4203387.588,125
628705.994,4204362.582,126
628727.292,4205307.577,127
629111.385,4206191.569,128
629855.074,4206984.558,129
630653.664,4207075.552,130
630870.066,4207868.542,131
630187.276,4207929.546,132
630138.585,4209178.534,133
629163.213,4211556.517,134
630394.572,4204515.569,135
627054.050,4213202.515,37
643007.132,4200888.461,138
642345.728,4202381.463,139
635487.739,4205825.516,140
634030.847,4205002.534,141
633945.452,4203692.542,142
632397.057,4203661.558,143
631110.866,4203661.569,144
629794.082,4203631.578,145
637810.353,4199729.521,146
635920.551,4201833.532,147
634488.053,4202808.541,148
642979.812,4181259.520,154
642208.613,4181533.531,155
641931.310,4182264.533,156
641373.513,4181838.543,157
640008.013,4182417.562,159
639547.712,4183057.566,160
639285.610,4183666.568,149
648865.505,4180466.431,162
646829.401,4182142.459,163
645354.197,4183819.478,164
643500.996,4185038.502,165
645314.600,4183209.480,166
643500.997,4184703.503,167
641525.898,4185404.529,168
639538.604,4185160.558,169
640318.895,4186989.541,170
638228.000,4186958.570,171
635673.706,4186867.606,173
634357.009,4186836.624,174
633326.811,4186836.639,175
632150.214,4186806.655,176
630894.518,4186775.665,177
628824.926,4186745.677,178
625459.938,4186288.700,179
625085.040,4185831.704,180
624569.941,4184215.715,181
628343.325,4188513.671,182
628748.721,4189549.663,183
628940.719,4190098.659,184
628322.022,4190159.662,185
628358.521,4190951.658,186
627691.025,4190677.663,187
631924.690,4193999.618,188
630522.602,4193207.632,189
629663.109,4192749.640,190
628837.116,4192292.648,191
627303.926,4191378.662,192
623765.246,4188117.701,193
628977.305,4197169.620,194
627492.918,4197139.630,195
625121.639,4197657.644,196
624021.249,4197870.650,197
622521.663,4197535.662,198
622326.566,4198754.657,199
622134.570,4199912.652,200
622305.270,4201558.643,201
622686.267,4202686.634,202
623472.658,4203570.624,203
622558.270,4204088.628,204
620970.290,4204210.639,205
619367.009,4203997.651,206
628669.393,4207349.563,207
627032.718,4207898.570,208
622945.350,4188757.703,209
623868.846,4189153.695,210
624463.243,4189945.687,211
624923.441,4191286.678,212
627489.914,4200095.614,213
620970.291,4204515.637,214
620884.895,4206313.629,215
622280.886,4208630.596,216
621445.794,4207898.610,217
620385.107,4207624.621,218
621284.207,4210215.587,219
618211.854,4211860.591,220
616431.869,4210001.623,221
618958.628,4208111.626,222
615450.476,4208325.649,223
622524.807,4213415.544,224
620177.831,4212196.573,225
618586.753,4212805.578,226
590536.046,4213750.818,227
621174.521,4212775.560,230
623853.689,4213080.539,231
624155.378,4211708.551,232
621299.511,4210977.579,234
622424.200,4211708.563,235
615517.475,4208172.650,236
612320.218,4208386.671,237
588070.229,4215427.824,238
620171.765,4219633.494,239
615395.617,4219328.528,240
641879.422,4208477.439,241
638636.359,4211799.435,242
635158.579,4212775.456,243
633384.675,4211434.485,244
631345.607,4214756.470,245
638861.894,4216493.387,246
635176.891,4214482.439,247
634110.107,4216189.432,248
632217.330,4218505.425,249
632122.820,4217042.440,250
629827.738,4216585.462,251
627462.465,4216463.479,252
631549.955,4236214.250,253
631351.850,4235086.262,254
631537.741,4233715.275,255
631385.336,4233014.283,256
636551.739,4235269.219,257
633326.947,4235391.244,258
632592.338,4233623.267,259
631909.629,4232099.288,260
631891.316,4230301.307,261
633180.599,4228411.316,262
632269.190,4226948.338,263
632046.678,4225150.359,264
631104.871,4223473.383,265
631016.463,4222285.396,266
631296.852,4221157.405,267
631699.140,4219724.417,268
629266.869,4220334.427,269
626871.192,4219755.449,270
624816.922,4221157.447,271
624347.516,4219023.473,272
605245.781,4236976.423,273
635564.101,4229569.285,275
634454.575,4225637.334,277
637508.648,4223229.332,278
634533.851,4222407.366,279
630760.532,4231733.301,280
630928.120,4230301.314,281
630391.619,4229417.327,282
629145.026,4228746.341,283
628928.615,4226857.362,284
628788.408,4225515.377,285
627569.205,4223108.409,286
626240.314,4222376.425,287
628919.548,4231855.310,288
627840.556,4231551.319,289
628172.744,4230209.332,290
626852.944,4228228.360,291
624969.353,4226887.386,292
624082.351,4224936.412,293
623780.544,4223016.434,294
623158.744,4221797.451,295
628739.735,4252643.112,296
627633.330,4250326.145,297
626420.228,4247888.178,298
624725.531,4246059.208,299
623753.230,4243560.237,300
622719.930,4241243.264,301
621945.729,4238439.291,302
623268.618,4237342.291,303
622421.218,4234873.316,304
622308.507,4232221.344,305
620622.901,4228137.399,306
628051.032,4269071.011,309
623344.909,4266572.082,310
623488.071,4259165.107,311
621997.664,4254776.160,312
619714.661,4248802.229,313
616992.762,4236793.335,315
616017.459,4232160.382,316
616483.772,4243895.291,317
616745.966,4238622.324,318
614182.585,4243133.314,319
611582.601,4238622.359,320
614325.782,4235208.361,321
614731.176,4233715.371,322
615267.669,4233075.376,323
607129.500,4235391.412,324
609135.119,4235300.392,325
611430.204,4235208.379,326
587744.022,4223991.729,327
594099.169,4214268.777,328
586698.624,4214177.860,329
629904.270,4272880.970,330
628910.534,4269162.998,331
628623.992,4264591.014,332
625633.876,4262152.056,333
628532.561,4259409.049,334
630623.441,4255721.063,335
628383.141,4253892.104,336
629187.820,4249229.141,337
628264.212,4245937.180,338
624527.424,4243072.235,339
624743.816,4240573.255,340
627682.085,4237250.264,341
629763.852,4233440.289,343
626301.279,4233288.310,344
626273.866,4231002.334,345
626270.854,4229112.354,346
624067.064,4227314.387,347
622043.271,4224875.425,348
619586.599,4225698.432,349
616736.730,4226277.443,350
614843.934,4222528.496,351
613332.138,4218718.549,352
610418.264,4216250.596,353
605187.838,4212988.682,354
601076.114,4214055.710,355
597549.489,4211556.774,356
592300.857,4212714.813,357
585644.020,4213141.891,358
581023.203,4212379.983,359
577182.688,4210734.067,360
575853.783,4209728.098,361
588499.934,4212561.852,362
585650.119,4216981.849,363
582745.308,4220456.872,364
582632.508,4218871.890,365
584113.914,4215091.899,366
579898.499,4214939.981,367
584702.115,4218840.848,368
575244.190,4230362.952,369
575783.691,4230209.940,370
584851.511,4230606.718,371
584357.710,4229752.739,372
584205.310,4227527.767,373
583318.308,4226034.803,374
582056.505,4225241.839,375
582553.307,4223717.843,376
580389.201,4221248.914,377
581096.303,4219694.913,378
576527.392,4229447.928,379
577770.995,4227801.913,380
577819.694,4224693.939,381
578688.396,4223717.928,382
579237.097,4221462.936,383
578980.996,4218597.967,384
578724.995,4215823.996,385
579730.799,4223900.903,386
581431.603,4227344.833,387
581285.303,4226156.847,388
578938.397,4226826.895,389
580322.201,4226582.865,390
578414.095,4224906.924,391
583095.807,4231459.752,392
581358.503,4228807.820,393
582788.006,4228563.789,394
586180.413,4231276.679,395
578139.796,4231063.876,396
585046.612,4228929.732,397
585040.512,4227527.747,398
586671.117,4226521.721,399
586393.816,4226247.731,401
584589.411,4226217.772,402
593855.373,4230087.598,403
588545.726,4231154.639,404
587356.916,4231276.650,405
594720.979,4226125.635,406
596418.697,4231093.561,408
594775.881,4228503.607,409
595559.186,4226460.623,410
595696.386,4225424.634,412
591672.954,4226704.659,413
597918.395,4215579.724,415
597976.295,4214847.732,417
595610.984,4221949.674,420
593355.467,4224845.664,421
591301.051,4225333.678,422
588518.227,4226674.691,425
583086.708,4223382.835,428
593818.768,4216585.753,433
591517.552,4216920.773,434
588570.031,4218017.789,436
579791.799,4220151.936,438
579782.699,4218932.947,440
578840.796,4220273.955,442
579925.899,4223016.907,443
579221.797,4219359.955,444
581364.603,4223534.871,445
637130.839,4235482.212,446
637249.637,4235208.214,447
636405.454,4238134.193,448
634442.452,4236854.221,449
630888.586,4243072.187,450
631199.482,4242462.191,451
630166.182,4240999.213,452
630699.570,4238988.229,453
631470.658,4236915.243,454
630662.957,4235818.260,455
625645.831,4206831.591,98
630562.167,4205460.562,136
631156.558,4206130.554,137
618934.348,4236519.325,308
618431.454,4238744.312,307
631497.385,4211860.498,33
624976.567,4211592.546,101
618262.262,4244148.275,314
597598.92,4216803.34,418
630298,4234283,342
627302,4187963,72
633465.55,4194204.52,112
628267,4185764,69
636554,4186941,172
647151,4185852,8
;647228.685,4185800.446,8   ; Head of Old River Barrier
;628261.030,4185709.686,69  ; Old R @ Tracy Barrier
;627386.230,4187812.680,72  ; Clifton Court Forebay Intake Gates
;636444.904,4186897.595,172 ; Grant Line Canal Barrier
;630306.353,4234233.277,342 ; Delta Cross-Channel Gates
;597747.695,4216432.716,418 ; SMSCG/RRDS Gates