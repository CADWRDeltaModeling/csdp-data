﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      51
627898.6,4185906.3,OBD
635780.8,4193802,MTB
638631.8,4186457.6,DGL
627377.4,4187715.2,ORI
627243.2,4188117.2,WCI
628084.5,4186853.4,GLC
629291.6,4192502.2,VCU
637754.4,4187026.5,GLE
628312.5,4185763.1,OAD
649126.1,4183436.8,MSD
653005.8,4171637.9,SJR
639164.7,4183509.3,SUR
639228.5,4183752.9,TPI
639778,4185041,PDC
647096.2,4185827.7,OH1
638981.8,4184006.2,SGA
639555,4185573,PCCU
643229,4184985,PDUP
639072,4185270,PCCD
642021.8,4186071.2,ORX
640088,4185530,OTWW
635798.2,4185059.9,TWA
636491.6,4185281.5,OLD
643723.1587,4185003.321,PCNB
643589.2414,4184870.011,PCSB
632927.2,4194823.6,VIC
643018.6,4187320.1,UNI
642184.4,4193313.5,MHO
634779.4549,4193764.353,MRX
649512,4179437,DVI
642052.7,4188617.1,MRU
645200.2,4181269.9,TPP
648060.2,4187435.7,SJD
625718.9,4194688.9,OH4
628839.5,4200455,MDM
630537,4183977,ORM
642469,4181997,TPPA
632231.1776,4182733.49,OAAD
633766.8116,4183139.204,ORFU
630172.109,4186906.468,GLW
637086,4184987,OTBD
626952,4187911.6,CLC
605075.1,4208474.7,ANH
625406.5,4203423.6,BAC
610598.8,4215917.6,EMM
624614.6,4207543.5,HLL
624476.9,4208582.2,HOL
615024.3,4212414.2,JER
575432.5,4209227.7,MRZ
646735.2,4199969.7,SJG
639210.2727,4181357.384,DAR
