﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      20
590134.7,4227040.1,BDL
625718.9,4194688.9,OH4
615196.3,4218095.3,TSL
636491.6,4185281.5,OLD
647096.2,4185827.7,OH1
630762.5,4257477,FPT
616676.6,4208098.2,DSJ
636454.1,4186988.1,GCT
628312.5,4185763.1,OAD
649126.1,4183436.8,MSD
575432.5,4209227.7,MRZ
646735.2,4199969.7,SJG
625222.5,4203213.9,OBI
629664.2,4235427.1,SDC
615024.3,4212414.2,JER
643575.2,4202944.9,RRI
629727.3,4233179.3,GSS
597451.6,4219938,NSL
605075.1,4208474.7,ANH
614797.6,4223035.8,SRV
