﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      91
647500.8,4192114.6,BDT
638631.8,4186457.6,DGL
626882.7,4186454,DMC
649512,4179437,DVI
636454.1,4186988.1,GCT
627753,4186838.8,GLC2
637754.4,4187026.5,GLE
642184.4,4193313.5,MHO
642052.7,4188617.1,MRU
635780.8,4193802,MTB
632905.7,4194776.6,MUP
628312.5,4185763.1,OAD
627898.6,4185906.3,OBD
628312.5,4185763.1,ODM
647096.2,4185827.7,OH1
625718.9,4194688.9,OH4
636491.6,4185281.5,OLD
630537,4183977,ORM
642021.8,4186071.2,ORX
639778,4185041,PDC
643229,4184985,PDUP
638981.8,4184006.2,SGA
648060.2,4187435.7,SJD
647576.1,4186166.1,SJL
639164.7,4183509.3,SUR
639228.5,4183752.9,TPS
639228.5,4183752.9,TPI
645200.2,4181269.9,TPP
635798.2,4185059.9,TWA
629291.6,4192502.2,VCU2
652957.8,4171293.8,VNS
647500.8,4192114.6,BDT
638631.8,4186457.6,DGL
626882.7,4186454,DMC
649512,4179437,DVI
636454.1,4186988.1,GCT
627753,4186838.8,GLC2
637754.4,4187026.5,GLE
642184.4,4193313.5,MHO
642052.7,4188617.1,MRU
635780.8,4193802,MTB
632905.7,4194776.6,MUP
628312.5,4185763.1,OAD
627898.6,4185906.3,OBD
628312.5,4185763.1,ODM
647096.2,4185827.7,OH1
625718.9,4194688.9,OH4
636491.6,4185281.5,OLD
630537,4183977,ORM
642021.8,4186071.2,ORX
639778,4185041,PDC
643229,4184985,PDUP
638981.8,4184006.2,SGA
648060.2,4187435.7,SJD
647576.1,4186166.1,SJL
639164.7,4183509.3,SUR
639228.5,4183752.9,TPS
639228.5,4183752.9,TPI
635798.2,4185059.9,TWA
629291.6,4192502.2,VCU2
652957.8,4171293.8,VNS
621783.2,4292647.4,VON
621783.2,4292647.4,VON
614797.6,4223035.8,SRV
614797.6,4223035.8,SRV
634300.2,4194175,MAB
627377.4,4187715.2,ORI
575432.5,4209227.7,MRZ
575432.5,4209227.7,MRZ
627243.2,4188117.2,WCI
627243.2,4188117.2,WCI
649126.1,4183436.8,MSD
649126.1,4183436.8,MSD
642289.3,4188756.4,MRMOW
642289.3,4188756.4,MRMOW
594757.5,4211123.3,MAL
605075.1,4208474.7,ANH
615105,4224350,RVB
615196.3,4218095.3,TSL
617515.3,4228186.2,RYF
608116.21,4215165.61,M13
619281.8,4227913.6,SXS
635762.3,4206110.6,TRN
616952.5,4212848.6,FAL
624652.3,4214658.4,OSJ
627377.4,4187715.2,ORI
624476.9,4208582.2,HOL
625222.5,4203213.9,OBI
615029,4212420.9,SJJ
646735.2,4199969.7,SJG
636598.9,4186932.5,GLAB
