﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      17
647500.8,4192114.6,BDT
638631.8,4186457.6,DGL
636598.9,4186932.5,GLAB
627753,4186838.8,GLC2
594757.5,4211123.3,MAL
628839.5,4200455,MDM
642184.4,4193313.5,MHO
642289.3,4188756.4,MRMOW
635780.8,4193802,MTB
632905.7,4194776.6,MUP
627898.6,4185906.3,OBD
639778,4185041,PDC
643229,4184985,PDUP
647576.1,4186166.1,SJL
639228.5,4183752.9,TPS
639228.5,4183752.9,TPI
645200.2,4181269.9,TPP
