﻿;HorizontalDatum:  UTMNAD83;HorizontalZone:   10;HorizontalUnits:  Meters;VerticalDatum:    NAVD88;VerticalUnits:    USSurveyFeet;Filetype:          landmark;NumElements:      20
632231.1776,4182733.49,OAAD
628084.5,4186853.4,GLC
637754.4,4187026.5,GLE
634300.2,4194175,MAB
642052.7,4188617.1,MRU
649126.1,4183436.8,MSD
628312.5,4185763.1,ODM
636491.6,4185281.5,OLD
627377.4,4187715.2,ORI
630537,4183977,ORM
642021.8,4186071.2,ORX
624652.3,4214658.4,OSJ
638981.8,4184006.2,SGA
648060.2,4187435.7,SJD
647576.1,4186166.1,SJL
646735.2,4199969.7,SJG
615029,4212420.9,SJJ
629291.6,4192502.2,VCU
652957.8,4171293.8,VNS
627243.2,4188117.2,WCI
