﻿;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      28
615180.4,4216618.4,SLTRM004
583348,4226330,SLSUS012
605228,4237166.9,SLBAR002
653005.8,4171637.9,RSAN112
643018.6,4187320.1,OLD_MID
636491.6,4185281.5,ROLD059
605075.1,4208474.7,RSAN007
631586.4,4219845,RSMKL008
626573,4213393.1,RSAN037
615105,4224350,RSAC101
580303.5,4226742.3,SLCBN002
619885.2,4204031,SLRCK005
625406.5,4203423.6,ROLD024
623513.4,4218211.2,RSAN032
623598.2,4238356.2,SSS
600858.7,4214644.1,RSAC081
629291.6,4192502.2,CHVCT000
615024.3,4212414.2,RSAN018
585550.4,4212803.2,RSAC064
626882.7,4186454,CHDMC006
647500.8,4192114.6,RSAN072
610598.8,4215917.6,RSAC092
590134.7,4227040.1,SLMZU011
626952,4187911.6,CHSWP003
643575.2,4202944.9,RSAN058
616676.6,4208098.2,SLDUT007
594757.5,4211123.3,RSAC075
597451.6,4219938,SLMZU025
