﻿;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      265
561701.6,4180706.7,aamc1
654346.1435,4277827,afo
584140.23,4160290.79,alam
550895.2,4186802.8,alk
588638.9,4144156,alv
588609.4,4144155.7,alvz
605075.1,4208474.7,anc
605075.1,4208474.7,anh
605075.1,4208474.7,anh2
640504,4269986,awb
625406.5,4203423.6,bac
590134.7,4227040.1,bdl
647500.8,4192114.6,bdt
636491.3,4235314.6,ben
576633.3,4211159,benbr
620980,4210523,bet
620996.1,4210486.7,bet2
629615.4,4207043.7,bir
605228,4237166.9,bks
595754.7,4226377.9,bll
612410.9,4210203.7,blp
582201.4519,4228997,bts
605282.66,4213133.12,c10
583902.55,4213517.57,c16
591743.04,4212444.61,c24
567940.8,4212900.6,carqb
614881,4234438,cbs
609500.3,4239525.4,ccs
603778.3506,4287183,ccy
628727.8,4189748.3,cis
626952,4187911.6,clc
600858.7,4214644.1,cll
542639,4199638.8,cm
618511,4244595,cm62
620970,4251599.2,cm66
623525.5,4259677.4,cm72
613995.8,4206152.6,cnt
602123.11,4213753.24,co5
597605.9,4211894.6,confl
586311.2,4146794.6,coy
594910,4142276.1,coycr
600859.1,4214643.6,cse
579678,4223160,cyg
624214.6,4197656.5,dbi
638631.8,4186457.6,dgl
630802.2,4234030.6,dlc
577868.3,4151149.6,dmb
626882.7,4186454,dmc
616676.6,4208098.2,dsj
577828.8,4151167.7,dum
578096,4151478.4,dumbr
649512,4179437,dvi
616657.3,4235072.2,dws
610598.8,4215917.6,emm
610598.8,4215917.6,emm2
616952.5,4212848.6,fal
616952.5,4212848.6,fal2
618521.7,4214201.8,fct
618582,4291614,few
579121.895,4214883,flt
584692.1,4227881.3,fmb
630762.5,4257477,fpt
615789.9,4290918.9,fre
623008.4,4211892.7,frk
619475.5,4208005.7,frp
636454.1,4186988.1,gct
629219.1,4233351.8,ges
586167.6,4143575.3,gl
636598.9,4186932.5,glab
628084.5,4186853.4,glc
627753,4186838.8,glc2
628084.6,4186841.5,glcgs
637754.4,4187026.5,gle
626989.2,4245160.4,gln
580533.214,4219949.694,god
582761,4218277.6,grizzb
624430.5,4221190.9,gsm
629727.3,4233179.3,gss
594479.1,4136908.3,guad
579253,4219416,gys
586986.9,4219943,gzb
584309.0232,4220037.891,gzl
582354,4221910,gzm
611430.5,4239220.3,has
623690.4,4187532.5,hbp
624614.6,4207543.5,hll
630093.3163,4208185.229,hlt
630737.3,4207200.2,hlt2
624476.9,4208582.2,hol
624476.9,4208582.2,hol2
624631.5,4203880,holm
593045.1,4214379.2,hon
623690.4,4187532.5,hro
585680,4231386,hsl
637297.2836,4270084,hst
582994.8199,4223547.67,hun
619734.2,4239063.4,hwb
577650.9,4223639,ibs
625220.4,4194097.8,idb
613977.7,4206196.5,inb
623050.7,4188795.5,ish
630173.3,4272187.3,ist
615024.3,4212414.2,jer
610819.69,4295934.45,klup
611458.99,4295736.72,knl
618409.8,4245456.2,lbtoe
616465,4243143,lct
616555,4239591,lcts
616465.4,4243142.6,lcut
617274,4243882,lhtn
617274,4243882,lhtse
615115,4233613,lib
616502.5,4242438.4,libc
614165.7,4242805.8,lir
623124,4259467.4,lis
623045.3,4262253.4,liw
614160.9,4243144.8,liy
631868.1,4217577.6,lps
608116.21,4215165.61,m13
634300.2,4194175,mab
594757.5,4211123.3,mal
565785.8,4213847.2,mare
566147.7,4159966.4,mateo
628839.5,4200455,mdm
628839.5,4200455,mdmzq
618522.3,4238860.6,mfv
670551,4263137,mhb
642184.4,4193313.5,mho
642165.8,4193399.5,mhr
616742.9,4232844.4,mir
630666.9,4231648.1,mkn
594844.5,4211136.4,mld
625274.8,4218552.5,mok
625274.8,4218552.5,mok2
585491.4,4149116.2,mow
642289.3,4188756.4,mrmow
642052.7,4188617.1,mru
634779.4549,4193764.353,mrx
575432.5,4209227.7,mrz
576774.9,4210025.7,mrz2
649126.1,4183436.8,msd
649126.1,4183436.8,msd2
597578.3032,4216762.676,msl
616742.4,4232792.7,mss
635780.8,4193802,mtb
599422.8,4051630.4,mtyc1
582570.3,4222664.5,mtz
632905.7,4194776.6,mup
560869,4246934.1,napr
630666.9,4231648.1,nmr
597451.6,4219938,nsl
597451.6,4219938,nsl2
581128.9,4152179.4,nw
628312.5,4185763.1,oad
627898.6,4185906.3,obd
625222.5,4203213.9,obi
628312.5,4185763.1,odm
647096.2,4185827.7,oh1
625718.9,4194688.9,oh4
636491.6,4185281.5,old
625738.9,4194696.3,orb
627355.1,4187787.9,orccf
627377.4,4187715.2,ori
630537,4183977,orm
625994.6,4209807.9,orq
625994.6,4209807.9,orq2
642021.8,4186071.2,orx
624652.3,4214658.4,osj
624652.3,4214658.4,osj2
585550.4,4212803.2,pct
580133.2256,4263389,pcw
639778,4185041,pdc
643229,4184985,pdup
531489.6,4232341.6,petr
590250.4,4142398,pond
627213.4,4213060.7,ppt
626573,4213393.1,pri
502341.4,4205260.6,pryc1
615325,4233252,psf
584266.1,4212463.8,ptchi
597238.3,4211183.7,pts
610695,4294664.3,rcs
548648.5,4198778.5,richb
552736,4198019.3,richm
638779.3,4206684.9,rindg
615252.9,4224292.9,riv
643575.2,4202944.9,rri
643575.2,4202944.9,rri2
621194.1,4204133.5,rsd
619885.2,4204031,rsl
569646.3,4151469.7,rtyc1
615105,4224350,rvb
588041.6,4215616.3,ryc
617515,4228186,rye
617515.3,4228186.2,ryf
616525.5,4230277.3,ryi
625540.70,4217496.70,sal
547485.2,4206082.9,scqc1
629664.2,4235427.1,sdc
610748.9,4216702.8,sdi
547094.8,4184503.1,sffpx
553143.4,4184169.8,sfp17
638981.8,4184006.2,sga
614250.8,4241943.7,sgg
550775.4,4196680.1,sham
641772,4204855,sjc
648060.2,4187435.7,sjd
646735.2,4199969.7,sjg
615029,4212420.9,sjj
647576.1,4186166.1,sjl
653005.8,4171637.9,sjr
586311.2,4146794.6,sm
632073.2,4231917.6,smr
632098.1,4231887.1,smr2
580303.5,4226742.3,snc
628119.1,4245666.2,snod
617644.9,4226137.5,soi
615180.4,4216618.4,sr3
629247.7,4247651,srh
614797.6,4223035.8,srv
623502,4218217,ssa
608608.2,4214765.6,ssi
623598.2,4238356.2,sss
617982,4243947,sstw
625441.04,4274267.15,ssw
626181,4255656,ssw2
631586.4,4219845,sti
639164.7,4183509.3,sur
622318.4,4234477.5,sus
624348.3,4243212.4,sut
629874.3,4233686.1,swe
619281.8,4227913.6,sxs
580045,4225811,tea
548699,4193884.8,tibc1
613974.4,4218374.1,tms
619009.8,4247207.4,toen
617130,4239083,toes
639228.5,4183752.9,tpi
645200.2,4181269.9,tpp
639228.5,4183752.9,tps
635762.3,4206110.6,trn
635762.3,4206110.6,trn2
626865,4186450,trp
615196.3,4218095.3,tsl
615192.5278,4218085.215,tss
635798.2,4185059.9,twa
616731,4217465,twi
612908.6,4237177.1,ucs
608463.8,4239164.3,ulc
643018.6,4187320.1,uni
629291.6,4192502.2,vcu
629291.6,4192502.2,vcu2
653005.8,4171637.9,ver
632927.2,4194823.6,vic
631822.4,4212328.2,vni
652957.8,4171293.8,vns
583348,4226330,vol
621783.2,4292647.4,von
621783.2,4292647.4,von2
648720,4224775,wbr
627243.2,4188117.2,wci
623426.6,4202761.2,wdcut
601759.47,4318532.21,wlk
610653.3539,4272076,wsd
618033.7,4281893.8,yby
