﻿;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      20
615180.4,4216618.4,SLTRM004
636491.6,4185281.5,ROLD059
605075.1,4208474.7,RSAN007
614797.6,4223035.8,RSAC101
625222.5,4203213.9,ROLD024
576774.9,4210025.7,RSAC054
646735.2,4199969.7,RSAN063
636454.1,4186988.1,CHGRL009
629727.3,4233179.3,Georg_SL
615029,4212420.9,RSAN018
625718.9,4194688.9,ROLD034
590134.7,4227040.1,SLMZU011
629664.2,4235427.1,RSAC128
630762.5,4257477,RSAC155
643575.2,4202944.9,RSAN058
616676.6,4208098.2,SLDUT007
628312.5,4185763.1,ROLD047
649126.1,4183436.8,RSAN087
647096.2,4185827.7,ROLD074
597451.6,4219938,SLMZU025
